module LightPattern3(clock,enable,greenLight, redLight);
	input clock, enable;
	output reg [0:7] greenLight, redLight;
	wire timer;
	
	reg [1:0]pattern; // remeber the flashing pattern.
	
	initial
	begin 
		pattern = 3'b0;
		greenLight = 8'b10010101;
		redLight = 8'b10101001;
	end
	
	PatternClock2 clk (timer, clock & enable, 1'b1);
	
	
	always @ (posedge timer or negedge enable) //ten seconds
	begin
		if(!enable)
		begin
			pattern <= 3'b0;
			greenLight <= 8'b10010101;
			redLight <= 8'b10101001;
		end
		else
		begin
			pattern <= pattern+1;
			case (pattern)
				3'b000:
				begin
					greenLight <= 8'b11001111;
					redLight <= 8'b11110011;
				end
				3'b001:
				begin
					greenLight <= 8'b01100000;
					redLight <= 8'b00001100;
				end
				3'b010:
				begin
					greenLight <= 8'b00111111;
					redLight <= 8'b11111100;
				end
				3'b011:
				begin
					greenLight <= 8'b11001111;
					redLight <= 8'b11110011;
				end
				3'b100:
				begin
					greenLight <= 8'b01010101;
					redLight <= 8'b10101010;
				end
				3'b101:
				begin
					greenLight <= 8'b10101010;
					redLight <= 8'b01010101;
				end
				3'b110:
				begin
					greenLight <= 8'b11001100;
					redLight <= 8'b00110011;
				end
				3'b111:
				begin
					greenLight <= 8'b00110011;
					redLight <= 8'b11001100;
				end
			endcase
		end
	end
endmodule 


module PatternClock3 (out, in, reset);
	input in, reset;
	output reg out;
	parameter freq = 12500000; //2;// 500000 units = 1/100th sec
	integer count;
	
	initial
	begin
		count = 0;
		out = 1'b0;
	end
	
	always @ (posedge in or negedge reset)
	begin
		if (~reset)
		begin
			count = 0;
			out = 1'b0;
		end
		else
		begin
			count = count + 1;
			if (count == freq / 2)
			begin
				out = ~out;
				count = 0;
			end
		end
	end
endmodule
